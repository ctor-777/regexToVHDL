
        library IEEE;
        use IEEE.std_logic_1164.all;

        entity something is
            port(
                som: in Character,
                thing: out std_logic
        );
        end entity;
        